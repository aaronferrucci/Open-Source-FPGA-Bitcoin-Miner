
bind fpgaminer_sys_tb test_program test_program_inst();

